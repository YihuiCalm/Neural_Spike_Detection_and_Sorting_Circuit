**.subckt inverter_tb
Vin Vin GND PULSE(0 5 0 0 0 5ns 10ns)
VDD VDD GND 5v
x1 Vout Vin inverter
**** begin user architecture code


.control
save all
tran 1ns 50ns
plot v(Vin) v(Vout)
.endc


 .lib /home/ubuntulab/IC/PDK/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=1

**** end user architecture code
**.ends

* expanding   symbol:  /media/sf_share/final_project/inverter.sym # of pins=2
* sym_path: /media/sf_share/final_project/inverter.sym
* sch_path: /media/sf_share/final_project/inverter.sch
.subckt inverter  vout vin
*.ipin vin
*.opin vout
XM3 vout vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 vout vin GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
